module xd(
    output [31:0] PCF,
    input [31:0] PCF_next,
    input CLK, RESET,
);

pc pc_inst( // TODO: AGREGAR stallF
    .PCF_curr(PCF),
    .PCF(PCF_next),
    .CLK(CLK),
    .RESET(RESET)
);

// pasamos el pc al adder para sumarle 4

adder pc_plus_4_inst(
    .Q(PCPlus4F),
    .A(PCF),
    .B(32'd4)
);


reg [31:0] instF;

ins_mem IMEM(
    .ins(instF),
    .address(PCF)
);

reg [31:0] insD, PCD, PCPlus4D;

IFID IFID_inst( // CORREGIR LOGICA STALLING y flushin walde matate:3
    .insD(insD),
    .PCD(PCD),
    .PCPlus4D(PCPlus4D),
    .flushD(flushD),
    .stallD(stallD),
    .CLK(CLK),
    .reset(RESET),
    .insF(instF),
    .PCPlus4F(PCPlus4F),
    .PCF(PCF)
);

reg [6:0] op;
reg [2:0] f3;
reg [6:0] f7;
reg [4:0] add_1, add_2, add_3;
reg [4:0] rs1D, rs2D, rdD;
reg [24:0] raw_imm;

decoder decoder_inst(
    .op(op),
    .f3(f3),
    .f7(f7),
    .add_1(add_1),
    .add_2(add_2),
    .add_3(add_3),
    .raw_imm(raw_imm), 
    .ins(insD)
);

wire [31:0] rd1, rd2, rdW;

reg_file reg_file_inst(
    .r_data_1(rd1),
    .r_data_2(rd2),
    .add_1(add_1),
    .add_2(add_2),
    .add_3(rdW),
    .write_data(resultW),
    .CLK(CLK),
    .REG_WRITE_W(regWriteW)
);

// ahora este neurotico duplica el a1(rs1D), a2(rs2D) y a3(rdD)

always @ (*) begin
    rs1D = add_1;
    rs2D = add_2;
    rdD = add_3;
end

reg regWriteD, memWriteD, jumpD, branchD, ALUSrcD;
reg [1:0] resultSrcD;
reg [2:0] immSrcD;
reg [3:0] ALUControlD;

control_unit control_unit_inst(
    .RES_SRC_D(resultSrcD),
    .REG_WRITE_D(regWriteD),
    .MEM_WRITE_D(memWriteD),
    .ALU_CONTROL_D(ALUControlD),
    .ALU_SRC_D(ALUSrcD),
    .IMM_SRC_D(immSrcD),
    .JUMP_D(jumpD),
    .BRANCH_D(branchD),
    .op(op),
    .f3(f3),
    .f7(f7)
);

reg [31:0] extImmD;
extender extender_inst(
    .imm(extImmD),
    .raw_imm(raw_imm),
    .immSrc(immSrcD)
);

// bueno ya extendimos ahora toca pasarle las cosas al IDEX osea que ya fue ya

reg [31:0] rd1E, rd2E, pcE, rs1E, rs2E, rdE, extImmE, PCPlus4E;
reg regWriteE, memWriteE, jumpE, branchE, ALUsrcE;
reg [3:0] ALUcontrolE;
reg [1:0] ResultSrcE;

IDEX IDEX_inst(
    .rd1E(rd1E), 
    .rd2E(rd2E), 
    .pcE(pcE), 
    .rs1E(rs1E), 
    .rs2E(rs2E), 
    .rdE(rdE), 
    .extImmE(extImmE), 
    .PCPlus4E(PC_plus_4E),
    .regWriteE(regWriteE),
    .memWriteE(memWriteE),
    .jumpE(jumpE),
    .branchE(branchE),
    .ALUsrcE(ALUsrcE),
    .ALUcontrolE(ALUcontrolE),
    .ResultSrcE(ResultSrcE),
    .rd1(rd1),
    .rd2(rd2),
    .pcD(PCD),
    .rs1D(rs1D),
    .rs2D(rs2D),
    .rdD(rdD),
    .extImmD(extImmD),
    .PC_plus_4D(PCPlus4D),
    .flushE(flushE),
    .regWriteD(regWriteD),
    .memWriteD(memWriteD),
    .jumpD(jumpD),
    .branchD(branchD),
    .ALUsrcD(ALUSrcD),
    .CLK(CLK),
    .reset(RESET),
    .ALUcontrolD(ALUControlD),
    .ResultSrcD(ResultSrcD)
);

// aqui vamos preparando el primer valor para el mux
reg [31:0] srcAE;

mux1_alu m1(
    .srcAE(srcAE),
    .rd1E(rd1E),
    .resultW(resultW),
    .aluResultM(aluResultM),
    .forwardAE(forwardAE),
);

// aqui el otro 
reg [31:0] mux2_out;

mux2_alu m2(
    .mux2_out(mux2_out),
    .rd2E(rd2E),
    .resultW(resultW),
    .aluResultM(aluResultM),
    .forwardBE(forwardBE),
);

// mux final para srcBE

wire [31:0] srcBE;
assign srcBE = ALUsrcE ? extImmE : mux2_out;

// add la, la, u time

wire zero;

alu alu_inst(
    .ALUResultE(aluResultE),
    .ZERO(zero),
    .src_A(srcAE),
    .src_B(srcBE),
    .ALUControlE(ALUcontrolE)
);

assign PCSrcE = jumpE || (zero && branchE);

// el adder ese para el pc

wire [31:0] PCTargetE;

adder adder_branch(
    .Q(PCTargetE),
    .A(pcE),
    .B(extImmE)
);

// ahora el EXMEM osea execute y memory

reg [31:0] rdM, aluResultM, writeDataM, PCPlus4M;
reg regWriteM, memWriteM;
reg [1:0] ResultSrcM;

EXMEM exmem_inst(
    .rdM(rdM),
    .aluResultM(aluResultM),
    .writeDataM(writeDataM),
    .PCPlus4M(PCPlus4M),
    .regWriteM(regWriteM),
    .memWriteM(memWriteM),
    .ResultSrcM(ResultSrcM),
    .regWriteE(regWriteE),
    .memWriteE(memWriteE),
    .CLK(CLK),
    .ResultSrcE(ResultSrcE),
    .aluResultE(aluResultE),
    .writeDataE(writeDataE),
    .PCPlus4E(PCPlus4E),
    .rdE(rdE)
);

// toca el data memory :3

reg [31:0] readDataM;

data_mem data_mem_inst(
    .r_data(readDataM),
    .write_data(writeDataM),
    .res_add(aluResultM),
    .MEM_WRITE(memWriteM),
    .CLK(CLK)
);

// ahora el MEMWB osea memory y write back

reg [31:0] readDataW, aluResultW, rdW, PCPlus4W;
reg regWriteW;
reg [1:0] ResultSrcW;

MEMWB MEMWB_inst(
    .readDataW(readDataW),
    .aluResultW(aluResultW),
    .rdW(rdW),
    .PC_plus_4W(PCPlus4W),
    .regWriteW(regWriteW),
    .ResultSrcW(ResultSrcW),
    .readDataM(readDataM),
    .aluResultM(aluResultM),
    .rdM(rdM),
    .PC_plus_4M(PCPlus4M),
    .regWriteM(regWriteM),
    .CLK(CLK),
    .ResultSrcM(ResultSrcM)
);

// finalmente el mux del write back

result_mux result_mux_inst(
    .resultW(resultW),
    .ALUResultM(aluResultW),
    .readDataW(readDataW),
    .PCPlus4W(PCPlus4W),
    .RES_SRC_W(ResultSrcW)
);

// el pc mux :3

pc_mux pc_mux_inst(
    .PC_next(PCF_next),
    .PCPlus4F(PCPlus4F),
    .PCTargetE(PCTargetE),
    .PCSrcE(PCSrcE)
);

// hazard unit :V

// :3333

// para forwardAE 
forwarding forwarding_inst(
    .forwardNE(forwardAE),
    .rsXE(rs1E),
    .rdM(rdM),
    .rdW(rdW),
    .regWriteM(regWriteM),
    .regWriteW(regWriteW)
);

// para forwardBE

forwarding forwarding_inst(
    .forwarNE(forwardAE),
    .rsXE(rs2E),
    .rdM(rdM),
    .rdW(rdW),
    .regWriteM(regWriteM),
    .regWriteW(regWriteW)
);

// stalling unit 7w7

wire lwStall, stallF, stallD, flushE;

stalling stalling_inst(
    .lwStall(lwStall),
    .stallF(stallF),
    .stallD(stallD),
    .flushE(flushE),
    .rs1D(rs1D),
    .rs2D(rs2D),
    .rdE(rdE),
);

flushing flushing_inst(
    .flushD(flushD),
    .flushE(flushE),
    .lwStall(lwStall),
    .PCSrcE(PCSrcE),
);
endmodule